package test_pkg;

	import uvm_pkg::*;

	`include "uvm_macros.svh"
`include "ahb_trans.sv"
`include "ahb_agent_config.sv"
`include "apb_agent_config.sv"
`include "env_config.sv"
`include "ahb_drv.sv"
`include "ahb_mon.sv"
`include "ahb_seqr.sv"
`include "ahb_agent.sv"
`include "ahb_agent_top.sv"
`include "ahb_seq.sv"

`include "apb_trans.sv"
`include "apb_drv.sv"
`include "apb_mon.sv"
`include "apb_seqr.sv"
`include "apb_seq.sv"
`include "apb_agent.sv"
`include "apb_agent_top.sv"

`include "virtual_seqr.sv"
`include "virtual_seqs.sv"
`include "scoreboard.sv"

`include "env.sv"


`include "test.sv"

endpackage